


module abc_dq0(clk, rstn, a, b, c, d, q, zero);

input wire [32:0] a;
input wire [32:0] b;
input wire [32:0] c;

endmodule